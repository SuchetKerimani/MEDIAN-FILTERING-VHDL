----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:53:09 03/23/2025 
-- Design Name: 
-- Module Name:    min_comp - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity min_comp is
    Port ( rst,clk : in  STD_LOGIC;
           A,B,C : in  STD_LOGIC_VECTOR (7 downto 0);
           MIN : OUT  STD_LOGIC_VECTOR (7 downto 0));
end min_comp;

architecture Behavioral of min_comp is
COMPONENT Eight_ip_dff is
    Port ( rst,clk : in  STD_LOGIC;
           d : in  STD_LOGIC_VECTOR (7 downto 0);
           q : out  STD_LOGIC_VECTOR (7 downto 0));
end COMPONENT;
 
component PE_min is 
    Port ( rst,clk : in  STD_LOGIC;
           A,B : in  STD_LOGIC_VECTOR (7 downto 0);
           min: out  STD_LOGIC_VECTOR (7 downto 0));
end  component;

signal MIN_1,Q_1:  STD_LOGIC_VECTOR (7 downto 0) ; 
begin
u1: PE_min port map (rst,clk,A,B,MIN_1);
u2: Eight_ip_dff port map (rst,clk,C,Q_1);
u3: PE_min port map (rst,clk,MIN_1,Q_1,MIN);
end Behavioral;

